--Instruction ROM loaded with UART test program with self test program and memory accesses


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom_7 is
    generic (
        WORDS : integer := 1024   -- 256 * 4B = 1 KB
    );
    port (
        clk     : in  std_logic;
--        rst_n   : in  std_logic;

        req    : in  std_logic;
        we     : in  std_logic;
        addr   : in  std_logic_vector(9 downto 0);  -- word address
        wdata  : in  std_logic_vector(31 downto 0);

        ready  : out std_logic;
        valid  : out std_logic;
        rdata  : out std_logic_vector(31 downto 0)
    );
end entity;

architecture rtl of rom_7 is

type mem_t is array (0 to WORDS-1) of std_logic_vector(31 downto 0);

constant ROM_INIT : mem_t := (



0=>  x"1fc21197",
1=>  x"80018193",
2=>  x"0fc11117",
3=>  x"ff810113",
4=>  x"00010433",
5=>  x"110000ef",
6=>  x"0000006f",
7=>  x"00000013",
8=>  x"00000013",
9=>  x"fe010113",
10=> x"00812e23",
11=> x"02010413",
12=> x"00050793",
13=> x"fef407a3",
14=> x"00000013",
15=> x"100127b7",
16=> x"0007a703",
17=> x"010007b7",
18=> x"00f777b3",
19=> x"fe0798e3",
20=> x"100127b7",
21=> x"fef44703",
22=> x"00e7a023",
23=> x"fef44703",
24=> x"100127b7",
25=> x"10076713",
26=> x"00e7a023",
27=> x"100127b7",
28=> x"fef44703",
29=> x"00e7a023",
30=> x"00000013",
31=> x"01c12403",
32=> x"02010113",
33=> x"00008067",
34=> x"fd010113",
35=> x"02112623",
36=> x"02812423",
37=> x"03010413",
38=> x"fca42e23",
39=> x"00700793",
40=> x"fef42623",
41=> x"0600006f",
42=> x"fec42783",
43=> x"00279793",
44=> x"fdc42703",
45=> x"00f757b3",
46=> x"00f7f793",
47=> x"fef42423",
48=> x"fe842703",
49=> x"00900793",
50=> x"00e7ec63",
51=> x"fe842783",
52=> x"0ff7f793",
53=> x"03078793",
54=> x"0ff7f793",
55=> x"0140006f",
56=> x"fe842783",
57=> x"0ff7f793",
58=> x"03778793",
59=> x"0ff7f793",
60=> x"00078513",
61=> x"f31ff0ef",
62=> x"fec42783",
63=> x"fff78793",
64=> x"fef42623",
65=> x"fec42783",
66=> x"fa07d0e3",
67=> x"00000013",
68=> x"00000013",
69=> x"02c12083",
70=> x"02812403",
71=> x"03010113",
72=> x"00008067",
73=> x"fc010113",
74=> x"02112e23",
75=> x"02812c23",
76=> x"04010413",
77=> x"100107b7",
78=> x"fef42023",
79=> x"fe042623",
80=> x"fe042423",
81=> x"05200513",
82=> x"eddff0ef",
83=> x"04900513",
84=> x"ed5ff0ef",
85=> x"05300513",
86=> x"ecdff0ef",
87=> x"04300513",
88=> x"ec5ff0ef",
89=> x"05600513",
90=> x"ebdff0ef",
91=> x"03300513",
92=> x"eb5ff0ef",
93=> x"03200513",
94=> x"eadff0ef",
95=> x"04900513",
96=> x"ea5ff0ef",
97=> x"00a00513",
98=> x"e9dff0ef",
99=> x"00d00513",
100=>x"e95ff0ef",
101=>x"04d00513",
102=>x"e8dff0ef",
103=>x"06500513",
104=>x"e85ff0ef",
105=>x"06d00513",
106=>x"e7dff0ef",
107=>x"06f00513",
108=>x"e75ff0ef",
109=>x"07200513",
110=>x"e6dff0ef",
111=>x"07900513",
112=>x"e65ff0ef",
113=>x"02000513",
114=>x"e5dff0ef",
115=>x"05400513",
116=>x"e55ff0ef",
117=>x"06500513",
118=>x"e4dff0ef",
119=>x"07300513",
120=>x"e45ff0ef",
121=>x"07400513",
122=>x"e3dff0ef",
123=>x"00a00513",
124=>x"e35ff0ef",
125=>x"00d00513",
126=>x"e2dff0ef",
127=>x"fec42783",
128=>x"00d79713",
129=>x"fec42783",
130=>x"0057d793",
131=>x"00f74733",
132=>x"a5a5a7b7",
133=>x"5a578793",
134=>x"00f747b3",
135=>x"fcf42e23",
136=>x"fe042223",
137=>x"1bc0006f",
138=>x"fe442703",
139=>x"040047b7",
140=>x"00f707b3",
141=>x"00279793",
142=>x"fcf42c23",
143=>x"fe442783",
144=>x"00279713",
145=>x"fdc42783",
146=>x"00f747b3",
147=>x"fe442703",
148=>x"00f747b3",
149=>x"fcf42a23",
150=>x"fe442783",
151=>x"00279793",
152=>x"fe042703",
153=>x"00f707b3",
154=>x"fd442703",
155=>x"00e7a023",
156=>x"fe442783",
157=>x"00279793",
158=>x"fe042703",
159=>x"00f707b3",
160=>x"0007a783",
161=>x"fcf42823",
162=>x"fd442703",
163=>x"fd042783",
164=>x"00f70863",
165=>x"fe842783",
166=>x"00178793",
167=>x"fef42423",
168=>x"00d00513",
169=>x"d81ff0ef",
170=>x"04900513",
171=>x"d79ff0ef",
172=>x"05400513",
173=>x"d71ff0ef",
174=>x"03a00513",
175=>x"d69ff0ef",
176=>x"fec42503",
177=>x"dc5ff0ef",
178=>x"02000513",
179=>x"d59ff0ef",
180=>x"04100513",
181=>x"d51ff0ef",
182=>x"04400513",
183=>x"d49ff0ef",
184=>x"04400513",
185=>x"d41ff0ef",
186=>x"05200513",
187=>x"d39ff0ef",
188=>x"03a00513",
189=>x"d31ff0ef",
190=>x"03000513",
191=>x"d29ff0ef",
192=>x"07800513",
193=>x"d21ff0ef",
194=>x"fd842503",
195=>x"d7dff0ef",
196=>x"02000513",
197=>x"d11ff0ef",
198=>x"03000513",
199=>x"d09ff0ef",
200=>x"07800513",
201=>x"d01ff0ef",
202=>x"fd442503",
203=>x"d5dff0ef",
204=>x"07c00513",
205=>x"cf1ff0ef",
206=>x"03000513",
207=>x"ce9ff0ef",
208=>x"07800513",
209=>x"ce1ff0ef",
210=>x"fd042503",
211=>x"d3dff0ef",
212=>x"02000513",
213=>x"cd1ff0ef",
214=>x"04500513",
215=>x"cc9ff0ef",
216=>x"05200513",
217=>x"cc1ff0ef",
218=>x"05200513",
219=>x"cb9ff0ef",
220=>x"03a00513",
221=>x"cb1ff0ef",
222=>x"fe842503",
223=>x"d0dff0ef",
224=>x"fe842783",
225=>x"00078e63",
226=>x"fe842783",
227=>x"0ff7f713",
228=>x"100117b7",
229=>x"0f076713",
230=>x"00e7a023",
231=>x"0140006f",
232=>x"100117b7",
233=>x"fe442703",
234=>x"00275713",
235=>x"00e7a023",
236=>x"fc042623",
237=>x"0100006f",
238=>x"fcc42783",
239=>x"00178793",
240=>x"fcf42623",
241=>x"fcc42703",
242=>x"0016e7b7",
243=>x"35f78793",
244=>x"fee7d4e3",
245=>x"fe442783",
246=>x"00178793",
247=>x"fef42223",
248=>x"fe442703",
249=>x"1ff00793",
250=>x"e4e7f0e3",
251=>x"fec42783",
252=>x"00178793",
253=>x"fef42623",
254=>x"e05ff06f",


    others => (others => '0')
);

signal mem : mem_t := ROM_INIT;

begin
    -- sempre pronta (single-cycle memory)
    ready <= '1';

    process(clk)
    begin
        if rising_edge(clk) then
            
                --rdata <= (others => '0');

                valid <= '0';

                if req = '1' then

                    if we = '1' then
                        mem(to_integer(unsigned(addr))) <= wdata;
                    end if;

                    -- lettura sincrona
                    rdata <= mem(to_integer(unsigned(addr)));
                    valid <= '1';
                end if;
            end if;
    end process;

end architecture;
