library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom_3 is
    generic (
        WORDS : integer := 1024   -- 256 * 4B = 1 KB
    );
    port (
        clk     : in  std_logic;
--        rst_n   : in  std_logic;

        req    : in  std_logic;
        we     : in  std_logic;
        addr   : in  std_logic_vector(9 downto 0);  -- word address
        wdata  : in  std_logic_vector(31 downto 0);

        ready  : out std_logic;
        valid  : out std_logic;
        rdata  : out std_logic_vector(31 downto 0)
    );
end entity;

architecture rtl of rom_3 is

type mem_t is array (0 to WORDS-1) of std_logic_vector(31 downto 0);

constant ROM_INIT : mem_t := (



0=>x"1fc21197",
1=>x"80018193",
2=>x"0fc11117",
3=>x"ff810113",
4=>x"00010433",
5=>x"010000ef",
6=>x"0000006f",
7=>x"00000013",
8=>x"00000013",
9=>x"10010337",
10=>x"00032783",
11=>x"fe010113",
12=>x"00112e23",
13=>x"00812c23",
14=>x"00912a23",
15=>x"01212823",
16=>x"01312623",
17=>x"01412423",
18=>x"01512223",
19=>x"00100713",
20=>x"00e7a023",
21=>x"00400713",
22=>x"00e7a223",
23=>x"00700713",
24=>x"00e7a423",
25=>x"00a00713",
26=>x"00e7a623",
27=>x"00d00713",
28=>x"00e7a823",
29=>x"01000713",
30=>x"00e7aa23",
31=>x"01300713",
32=>x"00e7ac23",
33=>x"01600713",
34=>x"00e7ae23",
35=>x"01900713",
36=>x"02e7a023",
37=>x"01c00713",
38=>x"02e7a223",
39=>x"01f00713",
40=>x"02e7a423",
41=>x"02200713",
42=>x"02e7a623",
43=>x"02500713",
44=>x"02e7a823",
45=>x"100108b7",
46=>x"02800713",
47=>x"02e7aa23",
48=>x"0048a803",
49=>x"02b00713",
50=>x"02e7ac23",
51=>x"02e00713",
52=>x"02e7ae23",
53=>x"0007a283",
54=>x"0047a683",
55=>x"0087af83",
56=>x"00c7af03",
57=>x"00d28733",
58=>x"0107ae83",
59=>x"01f70733",
60=>x"0147ae03",
61=>x"01e70733",
62=>x"0187a503",
63=>x"01d70733",
64=>x"01c7a583",
65=>x"01c70733",
66=>x"0207a483",
67=>x"00a70733",
68=>x"0247a383",
69=>x"00b70733",
70=>x"0287a083",
71=>x"00970733",
72=>x"02c7a403",
73=>x"00770733",
74=>x"0307a603",
75=>x"00170733",
76=>x"0347a903",
77=>x"00870733",
78=>x"0387a983",
79=>x"00c70733",
80=>x"03c7aa03",
81=>x"01270733",
82=>x"0007aa83",
83=>x"01370733",
84=>x"01470733",
85=>x"00ea8ab3",
86=>x"0157a023",
87=>x"0047aa83",
88=>x"0092c2b3",
89=>x"00169693",
90=>x"00ea84b3",
91=>x"0097a223",
92=>x"0087a483",
93=>x"0056c6b3",
94=>x"002f9f93",
95=>x"00e482b3",
96=>x"0057a423",
97=>x"00c7a283",
98=>x"01f6c6b3",
99=>x"003f1f13",
100=>x"00e28fb3",
101=>x"01f7a623",
102=>x"0107af83",
103=>x"01e6c6b3",
104=>x"004e9e93",
105=>x"00ef8f33",
106=>x"01e7a823",
107=>x"0147af03",
108=>x"01d6c6b3",
109=>x"005e1e13",
110=>x"00ef0eb3",
111=>x"01d7aa23",
112=>x"0187ae83",
113=>x"01c6c6b3",
114=>x"00651513",
115=>x"00ee8e33",
116=>x"01c7ac23",
117=>x"01c7ae03",
118=>x"00a6c6b3",
119=>x"00759593",
120=>x"00ee0533",
121=>x"00a7ae23",
122=>x"0207a503",
123=>x"00b6c6b3",
124=>x"00139393",
125=>x"00e505b3",
126=>x"02b7a023",
127=>x"0247a583",
128=>x"00d3c3b3",
129=>x"00209093",
130=>x"00e586b3",
131=>x"02d7a223",
132=>x"0287a683",
133=>x"0070c0b3",
134=>x"00341413",
135=>x"00e686b3",
136=>x"02d7a423",
137=>x"02c7a683",
138=>x"00144433",
139=>x"00461613",
140=>x"00e686b3",
141=>x"02d7a623",
142=>x"0307a683",
143=>x"00864633",
144=>x"00591913",
145=>x"00e686b3",
146=>x"02d7a823",
147=>x"0347a683",
148=>x"00c94933",
149=>x"00699993",
150=>x"00e686b3",
151=>x"02d7aa23",
152=>x"0387a603",
153=>x"0129c9b3",
154=>x"007a1693",
155=>x"00e60633",
156=>x"02c7ac23",
157=>x"03c7a603",
158=>x"0136c6b3",
159=>x"00e6c6b3",
160=>x"00e60733",
161=>x"02e7ae23",
162=>x"002dc7b7",
163=>x"00d82023",
164=>x"6bf78793",
165=>x"00000013",
166=>x"00078713",
167=>x"fff78793",
168=>x"fe071ae3",
169=>x"00032783",
170=>x"0048a803",
171=>x"e29ff06f",

    others => (others => '0')
);

signal mem : mem_t := ROM_INIT;

begin
    -- sempre pronta (single-cycle memory)
    ready <= '1';

    process(clk)
    begin
        if rising_edge(clk) then
            
                --rdata <= (others => '0');

                valid <= '0';

                if req = '1' then

                    if we = '1' then
                        mem(to_integer(unsigned(addr))) <= wdata;
                    end if;

                    -- lettura sincrona
                    rdata <= mem(to_integer(unsigned(addr)));
                    valid <= '1';
                end if;
            end if;
    end process;

end architecture;
